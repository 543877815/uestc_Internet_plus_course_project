`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/11/12 17:06:18
// Design Name: 
// Module Name: INSTMEM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module INSTMEM(Addr, Inst);
    input [31:0] Addr;
    output [31:0] Inst;
    wire [31:0] Rom [31:0];
    //��ͨCPU
//    assign Rom[5'h00] = 32'b100011_00000_00001_00000_000000_01100;//ȡ��������$1=3
//    assign Rom[5'h01] = 32'b100011_00000_00010_00000_000000_01000;//ȡ��������$2=2
//    assign Rom[5'h02] = 32'b000000_00001_00010_00011_000001_00000;//$3=$1+$2=5
//    assign Rom[5'h03] = 32'b000000_00001_00010_00100_000001_00010;//$4=$1-$2=1
//    assign Rom[5'h04] = 32'b000000_00011_00010_00101_000001_00100;//$5=$2&$3=0
//    assign Rom[5'h05] = 32'b000000_00011_00010_00110_000001_00101;//$6=$2|$3=7  
//    assign Rom[5'h06] = 32'b001100_00011_00111_0000000000000010;//$7=$3&2=0
//    assign Rom[5'h07] = 32'b001101_00011_01000_0000000000000010;//$8=$3|2=7
//    assign Rom[5'h08] = 32'b001000_00110_01001_0000000000000010;//$9=$6+2=9
//    assign Rom[5'h09] = 32'b100011_01001_01010_0000000000001000;//ȡ��������$10=$9+1000=100.01=4
//    assign Rom[5'h0A] = 32'b000100_00110_01000_0000000000000001;//$6��$8�������ת������ڶ���
//    assign Rom[5'h0B] = 32'b100011_00000_01011_00000_000000_00100;//ȡ��������$11=1
//    assign Rom[5'h0C] = 32'b100011_00000_01100_00000_000000_00100;//ȡ��������$12=1
//    assign Rom[5'h0D] = 32'b000101_00010_00001_0000000000000001;//$1��$2���������ת������ڶ���
//    assign Rom[5'h0E] = 32'b100011_00000_01101_00000_000000_00100;//ȡ��������$13=1
//    assign Rom[5'h0F] = 32'b100011_00000_01110_00000_000000_00100;//ȡ��������$14=1
//    assign Rom[5'h10] = 32'b000010_00000_00000_00000_000000_01110;//��ת�������ڶ���ָ��;
    
    //д����ǰ������
    assign Rom[5'h00] = 32'b100011_00000_00001_00000_000000_00100;//ȡ��������$1=1
    assign Rom[5'h01] = 32'b100011_00000_00010_00000_000000_01000;//ȡ��������$2=2
    assign Rom[5'h02] = 32'b100011_00000_00011_00000_000000_01100;//ȡ��������$3=3
    assign Rom[5'h03] = 32'b100011_00000_00100_00000_000000_10000;//ȡ��������$4=4
    //�ڲ�ǰ��
    assign Rom[5'h04] = 32'b001000_00001_00010_0000000000000010;//addi $2,$1,2; $2 = $1 + 2 = 3 
    assign Rom[5'h05] = 32'b000000_00010_00100_00011_000001_00100;//and $3,$4,$2; $3 = $4 & $2 = 4 & 3 = 0
    assign Rom[5'h06] = 32'b100011_00010_01000_0000000000011100;//lw $8, 7($2); $8 = 7
    assign Rom[5'h07] = 32'b001101_00010_00110_0000000000000100;//ori $6,$2,20; $6 = $2 | 4 = 3 | 4 = 7
    assign Rom[5'h08] = 32'b000000_00100_00010_00101_000001_00000;//add $5, $4, $2; $5 = $2 + $4 = 7
    //Lwָ�������ð��
    assign Rom[5'h09] = 32'b100011_00000_01100_00000_000000_10000;//ȡ��������$12=4
    assign Rom[5'h0A] = 32'b001000_01100_01011_0000000000000001;//addi $11, $12, 1; $11 = $12 + 1 = 5;
    assign Rom[5'h0B] = 32'b001100_01100_01110_0000000000000010;//andi $14, $12 , 2; $14 = $12 & 2 = 0;
    
//    assign Rom[5'h12] = 32'hXXXXXXXX;
//    assign Rom[5'h14] = 32'hXXXXXXXX;
//    assign Rom[5'h15] = 32'hXXXXXXXX;
//    assign Rom[5'h16] = 32'hXXXXXXXX;
//    assign Rom[5'h17] = 32'hXXXXXXXX;
//    assign Rom[5'h18] = 32'hXXXXXXXX;
//    assign Rom[5'h19] = 32'hXXXXXXXX;
//    assign Rom[5'h1A] = 32'hXXXXXXXX;
//    assign Rom[5'h1B] = 32'hXXXXXXXX;
//    assign Rom[5'h1C] = 32'hXXXXXXXX;
//    assign Rom[5'h1D] = 32'hXXXXXXXX;
//    assign Rom[5'h1E] = 32'hXXXXXXXX;
//    assign Rom[5'h1F] = 32'hXXXXXXXX;
    
    assign Inst = Rom [Addr[6:2]];
endmodule
